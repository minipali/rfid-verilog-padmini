`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: toptest
// Aditional comments:
// Simulates query command. 
//next to be simulated- ack
//////////////////////////////////////////////////////////////////////////////////
module toptest();

      // Regular IO
  // Oscillator input, master reset, demodulator input
  reg  reset, clk, demodin;

  // Modulator output
  wire modout;
  
  ///
  wire pll_enable;
  wire [3:0] freq_channel;
  wire rforbase;
  wire [12:0] commandparsed;
  //// sampsens
  wire adc_sample;
  wire [2:0] sensorcode;

  // Functionality control
  reg use_q, comm_enable;
  wire tx_enable;

  wire epc_data_ready;
  wire [15:0] writedataout;

  // Debugging IO
  wire  debug_clk;
  wire debug_out;
  
  /*registers storing the commands, samples from the 2MHz clock*/
   
  //reg [1909:0] bitquery; //Q = 1 query command
  reg [1800:0] bitquery;
  reg [430:0] bitqueryrep;
  reg [1582:0] bitack;
  reg [1704:0] bittrns;
  reg [2158:0] bitsamp;
  ///// some reead sample data code
  wire morb_trans;
  wire [7:0] sensor_time_stamp;
  wire [7:0] bf_dur;
  //crc5
  wire crc5invalid, crc16invalid;
  wire bitout;
  
  wire calibration_control;
  
  wire [15:0] counter;
  reg counterenb;
  wire overflow;
  reg counterreset;
  
  wire [2:0] sel_target;
  wire [2:0] sel_action;
  wire [7:0] sel_ptr;
  //wire [7:0] sel_masklen;
  wire [15:0] mask;
  wire [1:0] readwritebank; 
  wire [7:0] readwriteptr;
  wire [7:0] readwords; 
  wire membitclk, packet_complete;
  reg membitsrc, memdatadone,sl_flag;
  
 

  
  
  
  
  parameter QUERYREP   = 13'b0000000000001;
  parameter ACK        = 13'b0000000000010;
  parameter QUERY      = 13'b0000000000100;
  parameter QUERYADJ   = 13'b0000000001000;
  parameter SELECT     = 13'b0000000010000;//4
  parameter NACK       = 13'b0000000100000;
  parameter REQRN      = 13'b0000001000000;//6
  parameter READ       = 13'b0000010000000;//7
  parameter WRITE      = 13'b0000100000000;//8
  parameter TRNS       = 13'b0001000000000;
  parameter SAMPSENS   = 13'b0010000000000;
  parameter SENSDATA   = 13'b0100000000000;//11
  parameter BFCONST    = 13'b1000000000000;
  
  
  reg [12:0] command;
  
           
    initial begin
        reset = 1;
        clk = 0;
        demodin = 1;
        use_q = 1;
        comm_enable = 1;
        
        
        counterenb = 1;
        counterreset = 1;                           
        command = QUERY;
        sl_flag = 0;
        
        #200
        reset = 0;
        counterreset = 0;
        
        #1600000
        
//        command = TRNS;
//        counterreset = 0;
//        command = QUERYREP;
//        counterreset = 0;
//        #1600000
        
        command = ACK;
        counterreset = 0;
        
//        command = SAMPSENS;
//        counterreset = 0;
        
        #2000000
        $finish;
    end
    
    always #200 clk = ~clk; //2.5MHz clock frequency, bit rate
    
    assign debug_clk = clk;


    initial begin
       //below query is for q=0
       bitquery = 1801'b1111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       //bitquery = 1862'b11111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000;
       
       //will only work for sl flag 0
       //bitquery = 1910'b11111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000;
       //q=0 but invalid crc5
       //bitquery = 1848'b111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       bitqueryrep = 431'b00000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       bitack = 1583'b00000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       bittrns =  1705'b1111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       bitsamp = 2159'b00000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;         
    end
    
    
    

    always@(posedge clk && !reset) begin
    //initial
        if(counter <= 16'd1800 && command == QUERY) begin
            bitquery <= bitquery >> 1;
            demodin = bitquery;  
            if(counter >= 1800) begin 
                counterreset <=1;
                command <= 13'd0;
            end    
        end
        else if(counter <= 16'd430 && command == QUERYREP) begin 
       
            bitqueryrep <= bitqueryrep >> 1;
            demodin = bitqueryrep; 
            if(counter >= 430) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd1582 && command == ACK) begin 
       
            bitack <= bitack >> 1;
            demodin = bitack; 
            if(counter >= 1582) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd1704 && command == TRNS) begin 
       
            bittrns <= bittrns >> 1;
            demodin = bittrns; 
            
            if(counter >= 1704) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd2158 && command == SAMPSENS) begin 
       
            bitsamp <= bitsamp >> 1;
            demodin = bitsamp; 
            
            if(counter >= 2158) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else demodin =1; 
        
       
    end
    
    counter16 c10(.clk(clk), .reset(counterreset), .enable(counterenb), .count(counter), .overflow(overflow));
    
    top tp(reset, clk, demodin, modout, // regular IO
           writedataout,  epc_data_ready,
           readwritebank, readwriteptr, readwords, membitclk, membitsrc, memdatadone,
           use_q, comm_enable, tx_enable,
           debug_clk, debug_out,
           commandparsed,
           ///transmit clock
           pll_enable, freq_channel, rforbase,
           ////from sample data
           adc_sample, sensorcode,
           morb_trans, sensor_time_stamp, bf_dur,
           //crc checks
           crc5invalid, crc16invalid, bitout,
           calibration_control,
           sel_target, sel_action, sel_ptr, mask,
           sl_flag, packet_complete);
           
//module top(reset, clk, demodin, modout, // regular IO
//           writedataout, epc_data_ready,
//           readwritebank, readwriteptr, readwords, membitclk, membitsrc, memdatadone, 
//           use_q, comm_enable, tx_enable,
//           debug_clk, debug_out,
//           rx_cmd,
//           ///transmit clock
//           pll_enable, freq_channel, rforbase,
//           ////from sample data
//           adc_sample, senscode,
//           /////
//           morb_trans, sensor_time_stamp, bf_dur,      
//           crc5invalid, crc16invalid, bitout,
//           calibration_control,
//           //select
//           sel_target, sel_action, sel_ptr, mask,
//           sl_flag, packet_complete);


endmodule
