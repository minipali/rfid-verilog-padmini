`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module MC_test();

  //inputs to the module
  reg  reset, clk, demodin;
  reg use_q, comm_enable;
  reg [3:0] debug_address;
  reg factory_reset;
  
  reg ADC_data_ready;//add
  reg [7:0] ADC_data;//add
  reg [15:0] mem_read_in;
  
  
  //outputs
  wire [15:0] mem_data_out;
  wire PC_B,WE,SE;
  wire [5:0] mem_address;
  wire [2:0] mem_sel;
  wire modout;   
  wire tx_enable;                  
  wire debug_out;  
  wire osc_enable_pll;                               
  wire pll_enable;
  wire [3:0] freq_channel; 
  wire rforbase;                           
  wire [2:0] senscode;                            
  wire morb_trans;
  wire [7:0] bf_dur;
  wire backscatter_const;
  wire bitout, calibration_control;                                          
  wire packet_complete;   
  //not ops yet
//  wire [12:0] rx_cmd; 
//  wire [2:0] sel_target, sel_action; 
//  wire [5:0] counter_EPC, temp, read_or_write, counter_s1,counter_s2;
//  wire [3:0]write_state, bit_counter;
//  wire [15:0] tx_out;
//  wire [7:0] sel_ptr;                             
//  wire [15:0] mask; 
//  wire membitsrc;
//  wire memdatadone;
//  wire epc_data_ready;
//  reg fakememdone;
//  reg fakebitsrc;
  
  
  //ONLY FOR SIMULATIONS
  /*registers storing the commands, samples from the 2MHz clock*/
   
  //reg [1909:0] bitquery; //Q = 1 query command
  reg [1800:0] bitquery;
  reg [430:0] bitqueryrep;
  reg [1582:0] bitack;
  reg [1198:0] bittrns;
  reg [1582:0] bitsamp;
  reg [4035:0] bitselect;
  reg [2987:0] bitreqrn;
  reg [4535:0] bitwrite;
  reg [4151:0] bitread;
  reg [3575:0] bitsensdata;
  
  
  wire [15:0] counter;
  reg counterenb;
  wire overflow;
  reg counterreset;
  
  reg [12:0] command;  
  parameter QUERYREP   = 13'b0000000000001;
  parameter ACK        = 13'b0000000000010;
  parameter QUERY      = 13'b0000000000100;
  parameter QUERYADJ   = 13'b0000000001000;
  parameter SELECT     = 13'b0000000010000;//4
  parameter NACK       = 13'b0000000100000;
  parameter REQRN      = 13'b0000001000000;//6
  parameter READ       = 13'b0000010000000;//7
  parameter WRITE      = 13'b0000100000000;//8
  parameter TRNS       = 13'b0001000000000;
  parameter SAMPSENS   = 13'b0010000000000;
  parameter SENSDATA   = 13'b0100000000000;//11
  parameter BFCONST    = 13'b1000000000000;
           
    initial begin
        reset = 1;
        factory_reset = 1;
        clk = 0;
        demodin = 1;
        use_q = 0;
        comm_enable = 1;
        debug_address = 4'd12;
        
        
        //take care of these later
        ADC_data_ready = 0;
        ADC_data = 8'd0;
        mem_read_in = 16'h0000;
        
        counterenb = 1;
        counterreset = 1;                           
        //command = QUERY;
        command = SELECT;
        
        #250
        factory_reset = 0;
        
        #400
        reset = 0;
        factory_reset = 0;
        counterreset = 0;
        
        #2000000
        
//        command = TRNS;
//        counterreset = 0;
//        command = QUERYREP;
//        counterreset = 0;
//        #1600000
        
        command = QUERY;
        counterreset = 0;
        
        #1600000
        command = ACK;
        counterreset = 0;
        mem_read_in = 16'h0000;
        
        #3000000
        command = REQRN;
        counterreset = 0;
        
        #2400000
        command = SAMPSENS;
        counterreset = 0;
        
        #729600
        ADC_data = 8'b00000100;
        
        #400
        ADC_data_ready = 1;
        
        //#305200
        #120000
        ADC_data_ready = 0;
        
        #2000000
        
        command = TRNS;
        counterreset = 0;
        
        #2000000
        command = WRITE;
        counterreset = 0;
        
        #2400000
        bitwrite = 4536'b000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000;
        command = WRITE;
        counterreset = 0;
        
        #2400000
        bitwrite = 4536'b000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000;
        command = WRITE;
        counterreset = 0;
        
        #2400000
        command = READ;
        counterreset = 0;
        mem_read_in = 16'h0000;
        
        #1828600
        mem_read_in = 16'hA00A;
        #400
        mem_read_in = 16'hF00F;
        
        #2000000
        command = BFCONST;
        counterreset = 0;
        
        #1000000
        command = SENSDATA;
        counterreset = 0;
        
        #2000000
        $finish;
    end
    
    always #200 clk = ~clk; //2.5MHz clock frequency, bit rate
    initial begin
       //below query is for q=0
       bitquery = 1801'b1111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       //bitquery = 1862'b11111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000;
       
       //will only work for sl flag 0
       //bitquery = 1910'b11111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000;
       //q=0 but invalid crc5
       //bitquery = 1848'b111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       
       //bitselect = 3772'b0000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000;
       bitselect = 4036'b1111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000;
       bitreqrn = 2988'b000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000;
       bitqueryrep = 431'b00000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       bitack = 1583'b00000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       bittrns =  1199'b00000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       bitsamp = 1583'b00000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
       bitwrite = 4536'b000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000;
       bitread = 4152'b000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000;
       bitsensdata = 3576'b000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000;        
    end
    
    
    

    always@(posedge clk && !reset) begin
    //initial
        if(counter <= 16'd1800 && command == QUERY) begin
            bitquery <= bitquery >> 1;
            demodin = bitquery;  
            if(counter >= 1800) begin 
                counterreset <=1;
                command <= 13'd0;
            end    
        end
        else if(counter <= 16'd430 && command == QUERYREP) begin 
       
            bitqueryrep <= bitqueryrep >> 1;
            demodin = bitqueryrep; 
            if(counter >= 430) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd1582 && command == ACK) begin 
       
            bitack <= bitack >> 1;
            demodin = bitack; 
            if(counter >= 1582) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd1198 && command == TRNS) begin 
       
            bittrns <= bittrns >> 1;
            demodin = bittrns; 
            
            if(counter >= 1198) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd1582 && command == SAMPSENS) begin 
       
            bitsamp <= bitsamp >> 1;
            demodin = bitsamp; 
            
            if(counter >= 1582) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd4035 && command == SELECT) begin 
       
            bitselect <= bitselect >> 1;
            demodin = bitselect; 
            
            if(counter >= 4035) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd2987 && command == REQRN) begin 
       
            bitreqrn <= bitreqrn >> 1;
            demodin = bitreqrn; 
            
            if(counter >= 2987) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd4535 && command == WRITE) begin 
       
            bitwrite <= bitwrite >> 1;
            demodin = bitwrite; 
            
            if(counter >= 4535) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd4151 && command == READ) begin 
       
            bitread <= bitread >> 1;
            demodin = bitread; 
            
            if(counter >= 4151) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd3575 && command == SENSDATA) begin 
       
            bitsensdata <= bitsensdata >> 1;
            demodin = bitsensdata; 
            
            if(counter >= 3575) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else if(counter <= 16'd3598 && command == BFCONST) begin 
       
            bitsensdata <= bitsensdata >> 1;
            demodin = bitsensdata; 
            
            if(counter >= 3598) begin 
                counterreset <=1;
                command <= 13'd0;
            end   
        end
        else demodin =1; 
        
       
    end
    
    counter16 c10(.clk(clk), .reset(counterreset), .enable(counterenb), .count(counter), .overflow(overflow));
    
    top_MC_mem top_with_memory_inst(
            //top and memory
           reset, clk, 
           
           //directly top
           demodin, 
           use_q,
           comm_enable,
           debug_address,
           
           //directly to memory
           factory_reset,
           ADC_data_ready, 
           ADC_data, 
           mem_read_in,
           
           //directly from memory
           mem_data_out,
           PC_B,WE,SE,
           mem_address,
           mem_sel,
           
           
           modout, // regular IO
           tx_enable,
           debug_out,
           osc_enable_pll,
           pll_enable,
           freq_channel,
           rforbase,
           senscode,
           morb_trans,
           bf_dur,
           backscatter_const,
           bitout, 
           calibration_control,
           packet_complete);
           
//module top_MC_mem(
//            //top and memory
//           input reset, clk, 
           
//           //directly top
//           input demodin, 
//           input use_q,
//           input comm_enable,
//           input [3:0] debug_address,
           
           
//           //directly to memory
//           input factory_reset,
//           input ADC_data_ready, 
//           input [7:0] ADC_data, 
//           input [15:0] mem_read_in,
           
//           //directly from memory
//           output wire [15:0] mem_data_out, //data is given to the memory
//           output wire PC_B,WE,SE,
//           output wire [5:0] mem_address,  //this will enable WL
//           output wire [2:0] mem_sel,
           
           
//           //directly from top
//           output wire modout, // regular IO
//           output wire tx_enable,
//           output wire debug_out,
//           output wire osc_enable_pll,
//           output wire pll_enable,
//           output wire [3:0] freq_channel,
//           output wire rforbase,
//           output wire [2:0] senscode,
//           output wire morb_trans,
//           output wire [7:0] bf_dur,
//           output wire backscatter_const,
//           output wire bitout, calibration_control,
//           output wire packet_complete);
endmodule
